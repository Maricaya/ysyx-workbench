module top(
    input a,
    input b,
    output f
);
    assign f = a ^ b; // f = a XOR b
endmodule
